Param Rathour (190070049), CMOS Inverter
.include CMOS.txt ; Includes Solar Cell Model
.param Wn = {30u} Wp = {60u} Len = {0.4u}
.param Vd = 2.6
* M drain gate source body cmos
Mn out in gnd gnd cmosn L=Len W=Wn AS={2*Wn*Len} PS={2*Wn+4*Len} AD={2*Wn*Len} PD={2*Wn+4*Len}
Mp out in Vdd Vdd cmosp L=Len W=Wp AS={2*Wp*Len} PS={2*Wp+4*Len} AD={2*Wp*Len} PD={2*Wp+4*Len}
C1 out gnd 0.05p
Vdd Vdd gnd Vd
Vin in gnd pulse(0 Vd 0 20p 20p 4n 8n)
* .dc Vin 0 Vd 0.01
.tran 1p 30n
.control
let Vddd = Vd
run
let mid = {Vddd*0.5}
meas tran tpr1 WHEN V(in) = mid CROSS = 2
meas tran tpr2 WHEN V(out) = mid CROSS = 2
let tpr = tpr2-tpr1
meas tran tpf1 WHEN V(in) = mid CROSS = 3
meas tran tpf2 WHEN V(out) = mid CROSS = 3
let tpf = tpf2-tpf1
let tp = (tpr + tpf)/2
print tpr tpf tp
plot V(out) V(in)
wrdata 443.txt V(out); V(in)
.endc
.end