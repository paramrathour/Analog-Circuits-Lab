Param Rathour (190070049), Switching behaviour
.include BC547a.txt ; Includes BJT
Q1 c b e bc547a
Rb in b 1k
Vin in gnd pulse(0 5 0 0 0 0.25u 0.5u)
Vdd dd gnd 5
Rc dd c 1k
Ve e gnd 0
.tran 0.1u 2u
.control
run
plot V(c) V(in)
let I_C = -I(Vdd)
let I_B = -I(Vin)
plot I_C, I_B
.endc
.end