Param Rathour (190070049), Zener Diode in Voltage Regulator Experiment

.include zener.txt ; Includes Diode Model
.include ua741.txt ; Includes OpAmp Model
.include bc547.txt ; Includes BJT Model
.include Diode_1N914.txt            ; Includes Diode Model

Vin in gnd sin(0 16.7 50 0 0) ; Source Vin
Vop op gnd dc 12 ; DC Source Vin
Von on gnd dc -12 ; DC Source Vin

D1 in outp 1N914                     ; Diode
D2 outn in 1N914                     ; Diode
D3 outn gnd 1N914                    ; Diode
D4 gnd outp 1N914                    ; Diode
RL outp outn 1k                       ; Resistor (assumed 1k)
CL outp outn 100u                       ; Capacitor

q1 outp b e bc547a
x1 mid1 mid2 op on b UA741
RS outp mid1 100            ; Resistor
R1 e mid2 3.4k              ; Resistor
R2 mid2 outn 5.6k             ; Resistor
xR outn mid1  DI_1N4734A          ; Diode
.tran 0.1m 100m                     ; Transient Analysis
.control
run
plot {V(e) - V(outn)} vs {V(outp) - V(outn)}
plot {V(e) - V(outn)} ;{V(outp) - V(outn)}
* plot I(VdR) vs {V(mid1) - V(mid3)}

.endc
.end