Param Rathour (190070049), schottky_bat85

.include schottky_bat85.cir ; Includes Diode Model
.include TL071.cir ; Includes OpAmp Model

Vdc dc1 gnd dc 0
Vin in gnd sin(0 0.5 100k 0 0) ; Source Vin
Vp1 p1 gnd dc 15
Vn1 n1 gnd dc -15
Vp2 p2 gnd dc 15
Vn2 n2 gnd dc -15
R1 in ni1 10k
R2 dc1 ni1 1k
X1 gnd ni1 p1 n1 duti TL071
RF ni1 duti 1k
X2 duti duto BAT85
RFB duto out 150k
CFB duto out 100p
X3 gnd duto p2 n2 out TL071
.dc Vdc 0 5 0.01            ; DC Analysis
.control
run
let pi = 3.1415
let k1 = 100p*(sqrt(1+1/(2*pi*100k*150k*100p)^2))
plot abs({k1* V(out)/V(duti)}) vs abs(V(duti))
let k2 = 2/((1.03e-10)*(1.602e-19))
let area = 1p
let Cdut = abs({k1* V(out)/V(duti)})
let C = Cdut / area
let VD1 = -2
let VD2 = -4
let y = 1/C^2
meas dc C1 FIND y WHEN V(duti) = VD1
meas dc C2 FIND y WHEN V(duti) = VD2
let slope = (C2 - C1) / (VD2 - VD1)
print slope
plot 1/C^2 vs V(duti)
let ND = k2/abs(slope)
print ND
let yintercept = 0.00505435
* meas dc yintercept FIND y WHEN V(duti) = -1e-3
let Vbi = yintercept*ND/k2
print Vbi
.endc
.end