Param Rathour (190070049), Lighted I/V characteristics of Solar Cell
.include Solar_Cell.txt ; Includes Solar Cell Model
R1 in out 0
X1 out gnd solar_cell IL_val = 8e-3          	; Solar Cell
Vdummy in gnd 0;
.dc R1 1 500 0.1            ; DC Analysis
.control
set temp = 65
run
let I_D = -I(Vdummy)
let V_D = V(out)
plot I_D vs V_D
wrdata 24.txt I_D vs V_D
.endc
.end