Param Rathour (190070049), I/V characteristics of Diode 1N914

.include Diode_1N914.txt ; Includes Diode Model
R1 in mid1 100              ; Resistor
R2 mid1 gnd 1k              ; Resistor
R3 mid3 gnd 100             ; Resistor
dR mid1 midR 1N914          ; Diode
VdR midR mid3 0             ; Dummy Voltage to measure I_d
Vin in gnd dc 0             ; DC source Vin
.dc Vin 0 5 0.01 temp 20 80 10
.control
run
let Vout = {V(mid1) - V(mid3)}
plot I(VdR) vs Vout

wrdata 112.txt I(VdR) vs Vout
.endc
.end