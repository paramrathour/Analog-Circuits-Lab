Param Rathour (190070049), I/V characteristics of Solar Cell

.include Solar_Cell.txt ; Includes Solar Cell Model

R1 in out 0
X1 out gnd solar_cell IL_val = 10e-3          	; Solar Cell
Vdummy in gnd 0;
.dc R1 1 500 0.1            ; DC Analysis
.control
run
let I_D = -I(Vdummy)
let V_D = V(out)
let Power = I_D*V_D
plot I_D vs V_D
plot Power vs V_D
let I_SC = minimum(I_D)
let V_OC = maximum(V_D)
let Pmax = minimum(Power)
let FF = Pmax / (I_SC*V_OC)
print I_SC V_OC FF
* print Pmax; -2.14771e-03
* i_sc = -9.87702e-03
* v_oc = 4.249854e-01
* ff = 5.116530e-01
.endc
.end