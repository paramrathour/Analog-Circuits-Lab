Param Rathour (190070049), Reverse Recovery Time of Schottky BAT85

.include schottky_BAT85.txt ; Includes Diode Model
R1 in mid1 100              ; Resistor
R2 mid1 gnd 1k              ; Resistor
R3 mid3 gnd 100             ; Resistor
xR mid1 midR BAT85          ; Diode
VdR midR mid3 0             ; Dummy Voltage to measure I_d
Vin in gnd pulse(-5 5 0 0 0 0.005m 0.01m)             ; Pulsed input Vin
.tran 0.001u 5.1u 4.99u            ; Transient Analysis
.control
run
plot I(VdR) ;vs {V(mid1) - V(mid3)}
meas trans Imin MIN I(Vdr)
* meas trans Izero MIN abs(I(Vdr))
* meas trans tdiff I(Vdr) VAL=0, I(Vdr) VAL = 0; RISE = 1
meas trans t2 WHEN I(Vdr) = -1e-5 RISE = 1
meas trans t1 WHEN I(Vdr) = Imin
print t2 - t1
.endc
.end