Param Rathour (190070049), I/V characteristics of BLUE LED

.include blue_5mm.txt   ; Includes Diode Model
R1 in mid1 100               ; Resistor
R2 mid1 gnd 1k               ; Resistor
R3 mid3 gnd 100               ; Resistor
DB mid1 midB BLUE           ; Diode
VdB midB mid3 0 ; Dummy Voltage to measure I_d
Vin in gnd dc 0 ; DC source Vin
.dc Vin 0 5 0.01             ; DC Analysis
.control
run
let Vout = V(mid1) - V(mid3)
let VD1 = 2
let VD2 = 2.5
meas dc ID1 FIND I(VdB) WHEN Vout = VD1
meas dc ID2 FIND I(VdB) WHEN Vout = VD2
let lnID1 = log(ID1)
let lnID2 = log(ID2)
let eta = (VD2 - VD1) / ((26/1000) * (lnID2 - lnID1))
print lnID2 - lnID1
print eta
plot log(abs(I(VdB))) vs Vout
* wrdata B.txt log(abs(I(VdB))) Vout
.endc
.end