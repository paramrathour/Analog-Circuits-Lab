Param Rathour (190070049), BJT Parameters in CB configuration
.include BC547.txt ; Includes BJT
Q1 e b c bc547a
R1 mid c 100
Ib gnd b 1m
V2 mid gnd 0
V1 e gnd 2
.dc V2 0 20 0.01          ; DC Analysis
.control
run
let I_E = -I(V2)
let V_BC = {V(c) - V(b)}
plot I_E vs V_BC
wrdata 12b1.txt I_E vs V_BC
.endc
.end