Param Rathour (190070049), RC Lowpass
* Elements
* For Input Voltage as sin Wave with amplitude = 1V and Frequency Range 1Hz - 10kHz
Vin in gnd dc 0 ac 1
R1 in out 10k
C1 out gnd 0.1u

.ac DEC 10 1 10k

* Analysis
.control
run

* Display
plot V(in) V(out)
.endc

.end