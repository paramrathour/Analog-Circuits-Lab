Param Rathour (190070049), RC Differentiator
* Elements
* For Pulse Width = 10ms and Simulation Time = 100ms
Vin in gnd pulse(0 5 0 0 0 0.5m 1m)
C1 in out 0.1u
R1 out gnd 10k
.tran 0.01m 6m

* Analysis
.control
run

* Display
plot V(in) V(out)
.endc

.end