Param Rathour (190070049), BJT Parameters in CE configuration
.include bc547a.txt ; Includes BJT
Q1 c b e bc547a
R1 mid b 470
Ib in2 mid 0.1
V2 in2 gnd 0
R2 in1 c 100
V1 in1 gnd 0
Ve e gnd 0
.dc V1 0 10 0.1 temp 25 55 10       ; DC Analysis
.control
run
let I_C = -I(V1)
let V_CE = {V(c) - V(e)}
meas dc IC FIND I_C WHEN V_CE = 3
plot IC
.endc
.end