Param Rathour (190070049), Diode-Based Bridge Rectifier

.include Diode_1N914.txt            ; Includes Diode Model
Vin in gnd sin(0 16.9705627 50 0 0) ; Source Vin

D1 in outp 1N914                     ; Diode
D2 outn in 1N914                     ; Diode
D3 outn gnd 1N914                    ; Diode
D4 gnd outp 1N914                    ; Diode
RL outp outn 1k                       ; Resistor (assumed 1k)

.tran 0.01m 0.12                     ; Transient Analysis
.control
run
plot V(in) {V(outp) - V(outn)}
plot {V(outp) - V(outn)} vs V(in)

hardcopy 21.eps V(in) {V(outp) - V(outn)}
hardcopy 22.eps {V(outp) - V(outn)} vs V(in)
.endc
.end