Param Rathour (190070049), Common-Source Amplifier
.model NXYAA5U nmos Level=1 Vto=1 KP=100u w=10u L=1u + Gamma=0 Phi=0.65 Lambda=0.01
M1 d g s gnd NXYAA5U
VDD Vdd gnd 12                                      ; Supply Voltage
Vdum Vdd Vdum 0
Vin in gnd sin(0 50m 1000 0 0)                      ; Input Voltage
R1 Vdd g 8.2k                                       ; Resistor
R2 g gnd 3.3k                                       ; Resistor
RD d Vdum 3.3k                                      ; Resistor
RS s gnd 1k                                         ; Resistor
C1 g in 10u                                         ; Capacitor
CS s gnd 100u                                       ; Capacitor
.tran 0.001m 10m                                    ; Transient Analysis
.control                                            ; Control Functions
run
plot v(d)
meas trans V01 avg v(d)                             ; Finds DC op value
meas trans V01pp max v(d)
meas trans Vinpp max v(in)
let Gain = (V01pp-V01) / Vinpp
print Gain
.endc
.end