Param Rathour (190070049), BJT Current Source.include bc557.txt                                  ; Includes BJT Model.include zener_B.txt                                ; Includes Zener 5.6V ModelQ1 c b e bc557ax1 b Vcc zener_BVCC Vcc gnd 12                                      ; Supply VoltageVDL c L 0                                           ; Dummy VoltageRE Vcc e 4.7k                                       ; ResistorRB b gnd 2.2k                                       ; ResistorRL L gnd 1k                                         ; Resistor.dc RL 1k 10k 1k                                    ; DC Analysis (sweep R_L).control                                            ; Control Functionsrunplot I(VDL) vs V(L).endc.end