Param Rathour (190070049), Wien-bridge oscillator.include IN914.txt           					: Includes Diode Model.include ua741.txt           					: Includes Op-amp ModelVCCp VCCp gnd 12             					: Supply VoltageVCCn VCCn gnd -12            					: Supply Voltagex1 Vp Vn VCCp VCCn Vo ua741  					: Operational AmplifierR1 gnd Vn 4.7k               					: ResistorR2 Vn Vo 10k                 					: ResistorRF1 Vo Vmid 4.7k             					: ResistorCF1 Vmid Vp 0.1u             					: CapacitorRF2 Vp gnd 4.7k              					: ResistorCF2 Vp gnd 0.1u              					: Capacitor.tran 0.01m 525m 500m        					: Transient Analysis.control                     					: Control Functionsrunmeas trans Vpeak max V(Vo)plot V(Vo).endc.end