Param Rathour (190070049), RC Integrator
* Elements
Vin in gnd pulse(0 5 0 0 0 5m 10m)
R1 in out 10k
C1 out gnd 0.1u
.tran 0.01m 50m

* Analysis
.control
run

* Display
plot V(in) V(out)
.endc

.end