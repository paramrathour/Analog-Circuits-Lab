Param Rathour (190070049), I_D - V_GS Characteristics of PMOS at V_DS = -5V
.include pmos.txt ; Includes Solar Cell Model
M1 d g gnd gnd ALD1107
VD mid gnd -5
Vdummy d mid 0
VG g gnd 0
.dc VG 0 -5 -0.01           ; DC Analysis
.control
run
let I_D = I(Vdummy)
let V_GS = V(g)
plot sqrt(I_D) vs V_GS
wrdata 221.txt I_D vs V_GS
.endc
.end